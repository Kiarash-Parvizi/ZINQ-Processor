package types is
    type time_array is array(natural range <>) of time;
end package;
